-- de faup gregoire & estano paul

library ieee;
use ieee.std_logic_1164.all;
configuration fifo_test of fifo_tb is
  for fifo_tb_arch
  
  for DUT : FIFO
    for fifo1 
      for seqI: SEQ use entity 
        work.SEQ(Moore);
        --work.SEQ(Mealy);
      end for;
    end for;
  end for;
end for;
end fifo_test;